package multiplier2_pkg is
    constant N_BITS : natural := 8;
end package multiplier2_pkg;
