package multiplier1_1_pkg is
    constant n_BITS : natural := 4;
end package multiplier1_1_pkg;
