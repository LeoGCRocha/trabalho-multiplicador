package multiplier2_pkg is
    constant n_BITS : natural := 8;
end package multiplier2_pkg;
