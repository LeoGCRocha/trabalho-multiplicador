package multiplier_pkg is
    constant n_BITS : natural := 8;
end package multiplier_pkg;
