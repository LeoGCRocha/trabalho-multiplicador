package multiplier_pkg is
    constant n_BITS : natural := 16;
end package multiplier_pkg;
