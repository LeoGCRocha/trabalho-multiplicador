-- library ieee;
-- use ieee.std_logic_1164.all;
-- use ieee.numeric_std.all;
-- 
-- entity multiplier is
--     generic (n:natural => 4);
--     port(a, b   : in    signed(n-1 downto 0);
--         
